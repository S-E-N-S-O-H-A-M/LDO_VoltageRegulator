.lib "sky130_fd_pr/models/sky130.lib.spice" tt
xm3 net-_m1-pad1_ net-_m1-pad1_ gnd gnd sky130_fd_pr__nfet_01v8 W=0.42u L=0.5u
xm7 net-_m6-pad3_ net-_m1-pad1_ gnd gnd sky130_fd_pr__nfet_01v8 W=0.42u L=0.5u
xm2 net-_m1-pad1_ net-_m1-pad2_ net-_m2-pad3_ net-_m1-pad1_ sky130_fd_pr__pfet_01v8 W=3u L=0.5u
xm6 net-_m1-pad1_ net-_m2-pad3_ net-_m6-pad3_ net-_m1-pad1_ sky130_fd_pr__pfet_01v8 W=3u L=0.5u
xm1 net-_m1-pad1_ net-_m1-pad2_ net-_m1-pad2_ net-_m1-pad1_ sky130_fd_pr__pfet_01v8 W=3u L=0.5u
xm8 net-_m1-pad1_ net-_m6-pad3_ net-_c1-pad1_ net-_m1-pad1_ sky130_fd_pr__pfet_01v8 W=3u L=0.5u
xm5 net-_m4-pad3_ net-_m1-pad1_ gnd gnd sky130_fd_pr__nfet_01v8 W=0.42u L=0.5u
r1  net-_m9-pad2_ net-_c1-pad1_ 60k
r2  gnd net-_m9-pad2_ 100k
c1  net-_c1-pad1_ gnd 50pf
v2  vref gnd 1.50v
v1  net-_u2-pad1_ gnd 2.55v
* u4  vref plot_v1
* u2  net-_u2-pad1_ net-_m1-pad1_ plot_i2
xm4 net-_m1-pad2_ vref net-_m4-pad3_ net-_m4-pad3_ sky130_fd_pr__nfet_01v8 W=0.42u L=0.5u
xm9 net-_m2-pad3_ net-_m9-pad2_ net-_m4-pad3_ net-_m4-pad3_ sky130_fd_pr__nfet_01v8 W=0.42u L=0.5u
* u3  net-_c1-pad1_ gnd plot_i2
v_u2 net-_u2-pad1_ net-_m1-pad1_ 0
v_u3 net-_c1-pad1_ gnd 0
.tran 0e-00 100e-09 0e-09

* Control Statements 
.control
run
plot i(v_u2) i(v_u3)
.endc
.end
